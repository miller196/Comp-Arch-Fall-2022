module RAM(Addr, Write, Read, In, Out);

input [31:0] Addr;
input Write, Read;
input [31:0] In;  
output reg [31:0] Out; 

reg [31:0] RAM0, RAM1, RAM2, RAM3, RAM4, RAM5, RAM6, RAM7, RAM8, RAM9;
reg [31:0] RAM10, RAM11, RAM12, RAM13, RAM14, RAM15, RAM16, RAM17, RAM18, RAM19;
reg [31:0] RAM20, RAM21, RAM22, RAM23, RAM24, RAM25, RAM26, RAM27, RAM28, RAM29;
reg [31:0] RAM30, RAM31, RAM32, RAM33, RAM34, RAM35, RAM36, RAM37, RAM38, RAM39;
reg [31:0] RAM40, RAM41, RAM42, RAM43, RAM44, RAM45, RAM46, RAM47, RAM48, RAM49;
reg [31:0] RAM50, RAM51, RAM52, RAM53, RAM54, RAM55, RAM56, RAM57, RAM58, RAM59;
reg [31:0] RAM60, RAM61, RAM62, RAM63, RAM64, RAM65, RAM66, RAM67, RAM68, RAM69;
reg [31:0] RAM70, RAM71, RAM72, RAM73, RAM74, RAM75, RAM76, RAM77, RAM78, RAM79;
reg [31:0] RAM80, RAM81, RAM82, RAM83, RAM84, RAM85, RAM86, RAM87, RAM88, RAM89;
reg [31:0] RAM90, RAM91, RAM92, RAM93, RAM94, RAM95, RAM96, RAM97, RAM98, RAM99;
reg [31:0] RAM100, RAM101, RAM102, RAM103, RAM104, RAM105, RAM106, RAM107, RAM108, RAM109;
reg [31:0] RAM110, RAM111, RAM112, RAM113, RAM114, RAM115, RAM116, RAM117, RAM118, RAM119;
reg [31:0] RAM120, RAM121, RAM122, RAM123, RAM124, RAM125, RAM126, RAM127, RAM128, RAM129;
reg [31:0] RAM130, RAM131, RAM132, RAM133, RAM134, RAM135, RAM136, RAM137, RAM138, RAM139;
reg [31:0] RAM140, RAM141, RAM142, RAM143, RAM144, RAM145, RAM146, RAM147, RAM148, RAM149;
reg [31:0] RAM150, RAM151, RAM152, RAM153, RAM154, RAM155, RAM156, RAM157, RAM158, RAM159;
reg [31:0] RAM160, RAM161, RAM162, RAM163, RAM164, RAM165, RAM166, RAM167, RAM168, RAM169;
reg [31:0] RAM170, RAM171, RAM172, RAM173, RAM174, RAM175, RAM176, RAM177, RAM178, RAM179;
reg [31:0] RAM180, RAM181, RAM182, RAM183, RAM184, RAM185, RAM186, RAM187, RAM188, RAM189;
reg [31:0] RAM190, RAM191, RAM192, RAM193, RAM194, RAM195, RAM196, RAM197, RAM198, RAM199;
reg [31:0] RAM200, RAM201, RAM202, RAM203, RAM204, RAM205, RAM206, RAM207, RAM208, RAM209;
reg [31:0] RAM210, RAM211, RAM212, RAM213, RAM214, RAM215, RAM216, RAM217, RAM218, RAM219;
reg [31:0] RAM220, RAM221, RAM222, RAM223, RAM224, RAM225, RAM226, RAM227, RAM228, RAM229;
reg [31:0] RAM230, RAM231, RAM232, RAM233, RAM234, RAM235, RAM236, RAM237, RAM238, RAM239;
reg [31:0] RAM240, RAM241, RAM242, RAM243, RAM244, RAM245, RAM246, RAM247, RAM248, RAM249;
reg [31:0] RAM250, RAM251, RAM252, RAM253, RAM254, RAM255;

always @(Write)
begin
	case(Addr)
	32'd0 : RAM0 <= In;
	32'd1 : RAM1 <= In;
	32'd2 : RAM2 <= In;
	32'd3 : RAM3 <= In;
	32'd4 : RAM4 <= In;
	32'd5 : RAM5 <= In;
	32'd6 : RAM6 <= In;
	32'd7 : RAM7 <= In;
	32'd8 : RAM8 <= In;
	32'd9 : RAM9 <= In;
	32'd10 : RAM10 <= In;
	32'd11 : RAM11 <= In;
	32'd12 : RAM12 <= In;
	32'd13 : RAM13 <= In;
	32'd14 : RAM14 <= In;
	32'd15 : RAM15 <= In;
	32'd16 : RAM16 <= In;
	32'd17 : RAM17 <= In;
	32'd18 : RAM18 <= In;
	32'd19 : RAM19 <= In;
	32'd20 : RAM20 <= In;
	32'd21 : RAM21 <= In;
	32'd22 : RAM22 <= In;
	32'd23 : RAM23 <= In;
	32'd24 : RAM24 <= In;
	32'd25 : RAM25 <= In;
	32'd26 : RAM26 <= In;
	32'd27 : RAM27 <= In;
	32'd28 : RAM28 <= In;
	32'd29 : RAM29 <= In;
	32'd30 : RAM30 <= In;
	32'd31 : RAM31 <= In;
	32'd32 : RAM32 <= In;
	32'd33 : RAM33 <= In;
	32'd34 : RAM34 <= In;
	32'd35 : RAM35 <= In;
	32'd36 : RAM36 <= In;
	32'd37 : RAM37 <= In;
	32'd38 : RAM38 <= In;
	32'd39 : RAM39 <= In;
	32'd40 : RAM40 <= In;
	32'd41 : RAM41 <= In;
	32'd42 : RAM42 <= In;
	32'd43 : RAM43 <= In;
	32'd44 : RAM44 <= In;
	32'd45 : RAM45 <= In;
	32'd46 : RAM46 <= In;
	32'd47 : RAM47 <= In;
	32'd48 : RAM48 <= In;
	32'd49 : RAM49 <= In;
	32'd50 : RAM50 <= In;
	32'd51 : RAM51 <= In;
	32'd52 : RAM52 <= In;
	32'd53 : RAM53 <= In;
	32'd54 : RAM54 <= In;
	32'd55 : RAM55 <= In;
	32'd56 : RAM56 <= In;
	32'd57 : RAM57 <= In;
	32'd58 : RAM58 <= In;
	32'd59 : RAM59 <= In;
	32'd60 : RAM60 <= In;
	32'd61 : RAM61 <= In;
	32'd62 : RAM62 <= In;
	32'd63 : RAM63 <= In;
	32'd64 : RAM64 <= In;
	32'd65 : RAM65 <= In;
	32'd66 : RAM66 <= In;
	32'd67 : RAM67 <= In;
	32'd68 : RAM68 <= In;
	32'd69 : RAM69 <= In;
	32'd70 : RAM70 <= In;
	32'd71 : RAM71 <= In;
	32'd72 : RAM72 <= In;
	32'd73 : RAM73 <= In;
	32'd74 : RAM74 <= In;
	32'd75 : RAM75 <= In;
	32'd76 : RAM76 <= In;
	32'd77 : RAM77 <= In;
	32'd78 : RAM78 <= In;
	32'd79 : RAM79 <= In;
	32'd80 : RAM80 <= In;
	32'd81 : RAM81 <= In;
	32'd82 : RAM82 <= In;
	32'd83 : RAM83 <= In;
	32'd84 : RAM84 <= In;
	32'd85 : RAM85 <= In;
	32'd86 : RAM86 <= In;
	32'd87 : RAM87 <= In;
	32'd88 : RAM88 <= In;
	32'd89 : RAM89 <= In;
	32'd90 : RAM90 <= In;
	32'd91 : RAM91 <= In;
	32'd92 : RAM92 <= In;
	32'd93 : RAM93 <= In;
	32'd94 : RAM94 <= In;
	32'd95 : RAM95 <= In;
	32'd96 : RAM96 <= In;
	32'd97 : RAM97 <= In;
	32'd98 : RAM98 <= In;
	32'd99 : RAM99 <= In;
	32'd100 : RAM100 <= In;
	32'd101 : RAM101 <= In;
	32'd102 : RAM102 <= In;
	32'd103 : RAM103 <= In;
	32'd104 : RAM104 <= In;
	32'd105 : RAM105 <= In;
	32'd106 : RAM106 <= In;
	32'd107 : RAM107 <= In;
	32'd108 : RAM108 <= In;
	32'd109 : RAM109 <= In;
	32'd110 : RAM110 <= In;
	32'd111 : RAM111 <= In;
	32'd112 : RAM112 <= In;
	32'd113 : RAM113 <= In;
	32'd114 : RAM114 <= In;
	32'd115 : RAM115 <= In;
	32'd116 : RAM116 <= In;
	32'd117 : RAM117 <= In;
	32'd118 : RAM118 <= In;
	32'd119 : RAM119 <= In;
	32'd120 : RAM120 <= In;
	32'd121 : RAM121 <= In;
	32'd122 : RAM122 <= In;
	32'd123 : RAM123 <= In;
	32'd124 : RAM124 <= In;
	32'd125 : RAM125 <= In;
	32'd126 : RAM126 <= In;
	32'd127 : RAM127 <= In;
	32'd128 : RAM128 <= In;
	32'd129 : RAM129 <= In;
	32'd130 : RAM130 <= In;
	32'd131 : RAM131 <= In;
	32'd132 : RAM132 <= In;
	32'd133 : RAM133 <= In;
	32'd134 : RAM134 <= In;
	32'd135 : RAM135 <= In;
	32'd136 : RAM136 <= In;
	32'd137 : RAM137 <= In;
	32'd138 : RAM138 <= In;
	32'd139 : RAM139 <= In;
	32'd140 : RAM140 <= In;
	32'd141 : RAM141 <= In;
	32'd142 : RAM142 <= In;
	32'd143 : RAM143 <= In;
	32'd144 : RAM144 <= In;
	32'd145 : RAM145 <= In;
	32'd146 : RAM146 <= In;
	32'd147 : RAM147 <= In;
	32'd148 : RAM148 <= In;
	32'd149 : RAM149 <= In;
	32'd150 : RAM150 <= In;
	32'd151 : RAM151 <= In;
	32'd152 : RAM152 <= In;
	32'd153 : RAM153 <= In;
	32'd154 : RAM154 <= In;
	32'd155 : RAM155 <= In;
	32'd156 : RAM156 <= In;
	32'd157 : RAM157 <= In;
	32'd158 : RAM158 <= In;
	32'd159 : RAM159 <= In;
	32'd160 : RAM160 <= In;
	32'd161 : RAM161 <= In;
	32'd162 : RAM162 <= In;
	32'd163 : RAM163 <= In;
	32'd164 : RAM164 <= In;
	32'd165 : RAM165 <= In;
	32'd166 : RAM166 <= In;
	32'd167 : RAM167 <= In;
	32'd168 : RAM168 <= In;
	32'd169 : RAM169 <= In;
	32'd170 : RAM170 <= In;
	32'd171 : RAM171 <= In;
	32'd172 : RAM172 <= In;
	32'd173 : RAM173 <= In;
	32'd174 : RAM174 <= In;
	32'd175 : RAM175 <= In;
	32'd176 : RAM176 <= In;
	32'd177 : RAM177 <= In;
	32'd178 : RAM178 <= In;
	32'd179 : RAM179 <= In;
	32'd180 : RAM180 <= In;
	32'd181 : RAM181 <= In;
	32'd182 : RAM182 <= In;
	32'd183 : RAM183 <= In;
	32'd184 : RAM184 <= In;
	32'd185 : RAM185 <= In;
	32'd186 : RAM186 <= In;
	32'd187 : RAM187 <= In;
	32'd188 : RAM188 <= In;
	32'd189 : RAM189 <= In;
	32'd190 : RAM190 <= In;
	32'd191 : RAM191 <= In;
	32'd192 : RAM192 <= In;
	32'd193 : RAM193 <= In;
	32'd194 : RAM194 <= In;
	32'd195 : RAM195 <= In;
	32'd196 : RAM196 <= In;
	32'd197 : RAM197 <= In;
	32'd198 : RAM198 <= In;
	32'd199 : RAM199 <= In;
	32'd200 : RAM200 <= In;
	32'd201 : RAM201 <= In;
	32'd202 : RAM202 <= In;
	32'd203 : RAM203 <= In;
	32'd204 : RAM204 <= In;
	32'd205 : RAM205 <= In;
	32'd206 : RAM206 <= In;
	32'd207 : RAM207 <= In;
	32'd208 : RAM208 <= In;
	32'd209 : RAM209 <= In;
	32'd210 : RAM210 <= In;
	32'd211 : RAM211 <= In;
	32'd212 : RAM212 <= In;
	32'd213 : RAM213 <= In;
	32'd214 : RAM214 <= In;
	32'd215 : RAM215 <= In;
	32'd216 : RAM216 <= In;
	32'd217 : RAM217 <= In;
	32'd218 : RAM218 <= In;
	32'd219 : RAM219 <= In;
	32'd220 : RAM220 <= In;
	32'd221 : RAM221 <= In;
	32'd222 : RAM222 <= In;
	32'd223 : RAM223 <= In;
	32'd224 : RAM224 <= In;
	32'd225 : RAM225 <= In;
	32'd226 : RAM226 <= In;
	32'd227 : RAM227 <= In;
	32'd228 : RAM228 <= In;
	32'd229 : RAM229 <= In;
	32'd230 : RAM230 <= In;
	32'd231 : RAM231 <= In;
	32'd232 : RAM232 <= In;
	32'd233 : RAM233 <= In;
	32'd234 : RAM234 <= In;
	32'd235 : RAM235 <= In;
	32'd236 : RAM236 <= In;
	32'd237 : RAM237 <= In;
	32'd238 : RAM238 <= In;
	32'd239 : RAM239 <= In;
	32'd240 : RAM240 <= In;
	32'd241 : RAM241 <= In;
	32'd242 : RAM242 <= In;
	32'd243 : RAM243 <= In;
	32'd244 : RAM244 <= In;
	32'd245 : RAM245 <= In;
	32'd246 : RAM246 <= In;
	32'd247 : RAM247 <= In;
	32'd248 : RAM248 <= In;
	32'd249 : RAM249 <= In;
	32'd250 : RAM250 <= In;
	32'd251 : RAM251 <= In;
	32'd252 : RAM252 <= In;
	32'd253 : RAM253 <= In;
	32'd254 : RAM254 <= In;
	32'd255 : RAM255 <= In;
	endcase
end

always @(Read)
begin
	case(Addr)
	32'd0:Out <= RAM0;
	32'd1:Out <= RAM1;
	32'd2:Out <= RAM2;
	32'd3:Out <= RAM3;
	32'd4:Out <= RAM4;
	32'd5:Out <= RAM5;
	32'd6:Out <= RAM6;
	32'd7:Out <= RAM7;
	32'd8:Out <= RAM8;
	32'd9:Out <= RAM9;
	32'd10:Out <= RAM10;
	32'd11:Out <= RAM11;
	32'd12:Out <= RAM12;
	32'd13:Out <= RAM13;
	32'd14:Out <= RAM14;
	32'd15:Out <= RAM15;
	32'd16:Out <= RAM16;
	32'd17:Out <= RAM17;
	32'd18:Out <= RAM18;
	32'd19:Out <= RAM19;
	32'd20:Out <= RAM20;
	32'd21:Out <= RAM21;
	32'd22:Out <= RAM22;
	32'd23:Out <= RAM23;
	32'd24:Out <= RAM24;
	32'd25:Out <= RAM25;
	32'd26:Out <= RAM26;
	32'd27:Out <= RAM27;
	32'd28:Out <= RAM28;
	32'd29:Out <= RAM29;
	32'd30:Out <= RAM30;
	32'd31:Out <= RAM31;
	32'd32:Out <= RAM32;
	32'd33:Out <= RAM33;
	32'd34:Out <= RAM34;
	32'd35:Out <= RAM35;
	32'd36:Out <= RAM36;
	32'd37:Out <= RAM37;
	32'd38:Out <= RAM38;
	32'd39:Out <= RAM39;
	32'd40:Out <= RAM40;
	32'd41:Out <= RAM41;
	32'd42:Out <= RAM42;
	32'd43:Out <= RAM43;
	32'd44:Out <= RAM44;
	32'd45:Out <= RAM45;
	32'd46:Out <= RAM46;
	32'd47:Out <= RAM47;
	32'd48:Out <= RAM48;
	32'd49:Out <= RAM49;
	32'd50:Out <= RAM50;
	32'd51:Out <= RAM51;
	32'd52:Out <= RAM52;
	32'd53:Out <= RAM53;
	32'd54:Out <= RAM54;
	32'd55:Out <= RAM55;
	32'd56:Out <= RAM56;
	32'd57:Out <= RAM57;
	32'd58:Out <= RAM58;
	32'd59:Out <= RAM59;
	32'd60:Out <= RAM60;
	32'd61:Out <= RAM61;
	32'd62:Out <= RAM62;
	32'd63:Out <= RAM63;
	32'd64:Out <= RAM64;
	32'd65:Out <= RAM65;
	32'd66:Out <= RAM66;
	32'd67:Out <= RAM67;
	32'd68:Out <= RAM68;
	32'd69:Out <= RAM69;
	32'd70:Out <= RAM70;
	32'd71:Out <= RAM71;
	32'd72:Out <= RAM72;
	32'd73:Out <= RAM73;
	32'd74:Out <= RAM74;
	32'd75:Out <= RAM75;
	32'd76:Out <= RAM76;
	32'd77:Out <= RAM77;
	32'd78:Out <= RAM78;
	32'd79:Out <= RAM79;
	32'd80:Out <= RAM80;
	32'd81:Out <= RAM81;
	32'd82:Out <= RAM82;
	32'd83:Out <= RAM83;
	32'd84:Out <= RAM84;
	32'd85:Out <= RAM85;
	32'd86:Out <= RAM86;
	32'd87:Out <= RAM87;
	32'd88:Out <= RAM88;
	32'd89:Out <= RAM89;
	32'd90:Out <= RAM90;
	32'd91:Out <= RAM91;
	32'd92:Out <= RAM92;
	32'd93:Out <= RAM93;
	32'd94:Out <= RAM94;
	32'd95:Out <= RAM95;
	32'd96:Out <= RAM96;
	32'd97:Out <= RAM97;
	32'd98:Out <= RAM98;
	32'd99:Out <= RAM99;
	32'd100:Out <= RAM100;
	32'd101:Out <= RAM101;
	32'd102:Out <= RAM102;
	32'd103:Out <= RAM103;
	32'd104:Out <= RAM104;
	32'd105:Out <= RAM105;
	32'd106:Out <= RAM106;
	32'd107:Out <= RAM107;
	32'd108:Out <= RAM108;
	32'd109:Out <= RAM109;
	32'd110:Out <= RAM110;
	32'd111:Out <= RAM111;
	32'd112:Out <= RAM112;
	32'd113:Out <= RAM113;
	32'd114:Out <= RAM114;
	32'd115:Out <= RAM115;
	32'd116:Out <= RAM116;
	32'd117:Out <= RAM117;
	32'd118:Out <= RAM118;
	32'd119:Out <= RAM119;
	32'd120:Out <= RAM120;
	32'd121:Out <= RAM121;
	32'd122:Out <= RAM122;
	32'd123:Out <= RAM123;
	32'd124:Out <= RAM124;
	32'd125:Out <= RAM125;
	32'd126:Out <= RAM126;
	32'd127:Out <= RAM127;
	32'd128:Out <= RAM128;
	32'd129:Out <= RAM129;
	32'd130:Out <= RAM130;
	32'd131:Out <= RAM131;
	32'd132:Out <= RAM132;
	32'd133:Out <= RAM133;
	32'd134:Out <= RAM134;
	32'd135:Out <= RAM135;
	32'd136:Out <= RAM136;
	32'd137:Out <= RAM137;
	32'd138:Out <= RAM138;
	32'd139:Out <= RAM139;
	32'd140:Out <= RAM140;
	32'd141:Out <= RAM141;
	32'd142:Out <= RAM142;
	32'd143:Out <= RAM143;
	32'd144:Out <= RAM144;
	32'd145:Out <= RAM145;
	32'd146:Out <= RAM146;
	32'd147:Out <= RAM147;
	32'd148:Out <= RAM148;
	32'd149:Out <= RAM149;
	32'd150:Out <= RAM150;
	32'd151:Out <= RAM151;
	32'd152:Out <= RAM152;
	32'd153:Out <= RAM153;
	32'd154:Out <= RAM154;
	32'd155:Out <= RAM155;
	32'd156:Out <= RAM156;
	32'd157:Out <= RAM157;
	32'd158:Out <= RAM158;
	32'd159:Out <= RAM159;
	32'd160:Out <= RAM160;
	32'd161:Out <= RAM161;
	32'd162:Out <= RAM162;
	32'd163:Out <= RAM163;
	32'd164:Out <= RAM164;
	32'd165:Out <= RAM165;
	32'd166:Out <= RAM166;
	32'd167:Out <= RAM167;
	32'd168:Out <= RAM168;
	32'd169:Out <= RAM169;
	32'd170:Out <= RAM170;
	32'd171:Out <= RAM171;
	32'd172:Out <= RAM172;
	32'd173:Out <= RAM173;
	32'd174:Out <= RAM174;
	32'd175:Out <= RAM175;
	32'd176:Out <= RAM176;
	32'd177:Out <= RAM177;
	32'd178:Out <= RAM178;
	32'd179:Out <= RAM179;
	32'd180:Out <= RAM180;
	32'd181:Out <= RAM181;
	32'd182:Out <= RAM182;
	32'd183:Out <= RAM183;
	32'd184:Out <= RAM184;
	32'd185:Out <= RAM185;
	32'd186:Out <= RAM186;
	32'd187:Out <= RAM187;
	32'd188:Out <= RAM188;
	32'd189:Out <= RAM189;
	32'd190:Out <= RAM190;
	32'd191:Out <= RAM191;
	32'd192:Out <= RAM192;
	32'd193:Out <= RAM193;
	32'd194:Out <= RAM194;
	32'd195:Out <= RAM195;
	32'd196:Out <= RAM196;
	32'd197:Out <= RAM197;
	32'd198:Out <= RAM198;
	32'd199:Out <= RAM199;
	32'd200:Out <= RAM200;
	32'd201:Out <= RAM201;
	32'd202:Out <= RAM202;
	32'd203:Out <= RAM203;
	32'd204:Out <= RAM204;
	32'd205:Out <= RAM205;
	32'd206:Out <= RAM206;
	32'd207:Out <= RAM207;
	32'd208:Out <= RAM208;
	32'd209:Out <= RAM209;
	32'd210:Out <= RAM210;
	32'd211:Out <= RAM211;
	32'd212:Out <= RAM212;
	32'd213:Out <= RAM213;
	32'd214:Out <= RAM214;
	32'd215:Out <= RAM215;
	32'd216:Out <= RAM216;
	32'd217:Out <= RAM217;
	32'd218:Out <= RAM218;
	32'd219:Out <= RAM219;
	32'd220:Out <= RAM220;
	32'd221:Out <= RAM221;
	32'd222:Out <= RAM222;
	32'd223:Out <= RAM223;
	32'd224:Out <= RAM224;
	32'd225:Out <= RAM225;
	32'd226:Out <= RAM226;
	32'd227:Out <= RAM227;
	32'd228:Out <= RAM228;
	32'd229:Out <= RAM229;
	32'd230:Out <= RAM230;
	32'd231:Out <= RAM231;
	32'd232:Out <= RAM232;
	32'd233:Out <= RAM233;
	32'd234:Out <= RAM234;
	32'd235:Out <= RAM235;
	32'd236:Out <= RAM236;
	32'd237:Out <= RAM237;
	32'd238:Out <= RAM238;
	32'd239:Out <= RAM239;
	32'd240:Out <= RAM240;
	32'd241:Out <= RAM241;
	32'd242:Out <= RAM242;
	32'd243:Out <= RAM243;
	32'd244:Out <= RAM244;
	32'd245:Out <= RAM245;
	32'd246:Out <= RAM246;
	32'd247:Out <= RAM247;
	32'd248:Out <= RAM248;
	32'd249:Out <= RAM249;
	32'd250:Out <= RAM250;
	32'd251:Out <= RAM251;
	32'd252:Out <= RAM252;
	32'd253:Out <= RAM253;
	32'd254:Out <= RAM254;
	32'd255:Out <= RAM255;
	endcase
end

endmodule