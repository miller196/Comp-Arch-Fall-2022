module Multiplex_TB();

reg [4:0] Signal;

reg [31:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31;
wire [31:0] Output;

Multiplex dut (R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31, Signal, Output);

initial begin
	Signal <= 5'b00000;
	R0 <= 32'b00000000000000000000000000000001;
	R1 <= 32'b00000000000000000000000000000010;
	R2 <= 32'b00000000000000000000000000000100;
	R3 <= 32'b00000000000000000000000000001000;
	R4 <= 32'b00000000000000000000000000010000;
	R5 <= 32'b00000000000000000000000000100000;
	R6 <= 32'b00000000000000000000000001000000;
	R7 <= 32'b00000000000000000000000010000000;
	R8 <= 32'b00000000000000000000000100000000;
	R9 <= 32'b00000000000000000000001000000000;
	R10 <= 32'b00000000000000000000010000000000;
	R11 <= 32'b00000000000000000000100000000000;
	R12 <= 32'b00000000000000000001000000000000;
	R13 <= 32'b00000000000000000010000000000000;
	R14 <= 32'b00000000000000000100000000000000;
	R15 <= 32'b00000000000000001000000000000000;
	R16 <= 32'b00000000000000010000000000000000;
	R17 <= 32'b00000000000000100000000000000000;
	R18 <= 32'b00000000000001000000000000000000;
	R19 <= 32'b00000000000010000000000000000000;
	R20 <= 32'b00000000000100000000000000000000;
	R21 <= 32'b00000000001000000000000000000000;
	R22 <= 32'b00000000010000000000000000000000;
	R23 <= 32'b00000000100000000000000000000000;
	R24 <= 32'b00000001000000000000000000000000;
	R25 <= 32'b00000010000000000000000000000000;
	R26 <= 32'b00000100000000000000000000000000;
	R27 <= 32'b00001000000000000000000000000000;
	R28 <= 32'b00010000000000000000000000000000;
	R29 <= 32'b00100000000000000000000000000000;
	R30 <= 32'b01000000000000000000000000000000;
	R31 <= 32'b10000000000000000000000000000000;
	#1000 $stop;
	
end

	
always begin

	#5 Signal <= Signal + 5'b1;
	#5;
end

endmodule